module uartRx(
    input var logic clock,
    output var logic busy
);
endmodule
