module ram(
    
);
endmodule
